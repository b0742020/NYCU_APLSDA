//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//////////////////////////////////Lab04 Exercise//////////////////////////////
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   
//                       Author     		  : Hong-Ming Wu
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : FSM.v
//   Module Name : FSM
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module FSM(
    //Input Ports
    input [3:0]KEY,
    input [2:0]SW,
    //Output Ports
    output reg [6:0]HEX0  // Result output valid
);

//==============================================//
//             Parameter and Integer            //
//==============================================//
// State declaration for FSM
// Example: parameter IDLE = 3'b000;
parameter IDLE = 3'b000;
parameter RUNNING = 3'b001;
parameter PAUSE = 3'b010;
parameter FINISH = 3'b100;


//==============================================//
//                 reg declaration              //
//==============================================//
reg[3:0]result_ff,result;
reg[1:0]input_ff;


//==============================================//
//             Current State Block              //
//==============================================//



//==============================================//
//              Next State Block                //
//==============================================//



//==============================================//
//             Base and Score Logic             //
//==============================================//
// Handle base runner movements and score calculation.
// Update bases and score depending on the action:
// Example: Walk, Hits (1H, 2H, 3H), Home Runs, etc.



//==============================================//
//                Output Block                  //
//==============================================//
// Decide when to set out_valid high, and output score_A, score_B, and result.



endmodule
